module com_cc_rx(
    input clk,
    
    input fire_rxd,

    input pin_rxd,
    output reg usb_rxd
);

    





endmodule