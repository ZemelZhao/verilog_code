module console_usb(
    input clk,
    input rst
);



endmodule