module console_core(
    input clk,
    input rst,

    
);


endmodule