module top(
    input clk,
    input rst_n,


);

    wire rst;


    assign rst = ~rst_n;







    







endmodule
