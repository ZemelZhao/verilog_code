module tb_mactx(
    input clk,
    input rst
);

    


endmodule