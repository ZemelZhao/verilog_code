module com(
    input clk,
    input rst,

    input fs_send,
    output fd_send,
    output fs_read,
    input fd_read,

    
);




    eth
    eth_dut(
        .clk(),
        .rst(),

        .
    );


endmodule