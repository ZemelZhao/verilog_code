module trgg_in(

);
