module gmii_tx_buffer(
    input clk,
    input rst_n,
    input eth_100m_en,
    input eth_10m_en,

    input gmii_txen,
    input [7:0] gmii_txd,
    output e_100_txen,
    output [7:0] e_100_txd
); 




endmodule