module trgg(
    input clk,
    input rst,

    input fs,
    output fd,

    input [0:39] trgg_cmd,

    output [0:1] pin_trgg
);

    

endmodule