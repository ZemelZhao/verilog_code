module tb_inout(
    input clk,
    input rst_n,

    input [1:0] cc,

    inout [1:0] sbu
);

    reg state, next_state;

    
    



endmodule