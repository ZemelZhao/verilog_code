module top(
    input clk_in_p,
    input clk_in_n,

    input rst_n,
    output fan_n,

    output [0:5] led_stat_n,
    output [0:5] led_comm_n
);

    wire clk_slow, clk_norm, clk_fast, clk_ulta;

    



endmodule