module console_usb_sub(
    input clk,
    input rst


);



endmodule