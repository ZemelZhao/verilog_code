module top(
    input clk,
    input rst_n
);
    wire rst = ~rst_n;





endmodule