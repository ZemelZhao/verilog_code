module console_usb_hq(
    input clk,
    input rst
);


endmodule