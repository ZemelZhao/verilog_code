module com_cc(
    input clk_ulta,
    input clk_fast,

    input fire_rxd,
    input fire_txd,
    output pin_send,

    input [3:0] usb_txd,
    output [3:0] pin_txd,

    input pin_rxd,
    output usb_rxd
);

















endmodule
